`timescale 1ns / 1ps
module value_ROM(
    input [5:0] some_value, //МОДУЛЬ ВОСПРИНИМАЕТ ЧИСЛО В ВОСЬМЕРИЧНОЙ СИСТЕМЕ СЧИСЛЕНИЯ!
    input en,
    input newframe,
    output [7:0] exit_value
);
////////////////////////////////////////////////////////// 
wire [2:0] f_eight;
wire [2:0] s_eignt;
reg [7:0] value;
//////////////////////////////////////////////////////////
assign f_eight = some_value[2:0];
assign s_eignt = some_value[5:3];
assign exit_value = value;
//////////////////////////////////////////////////////////
always @(posedge newframe) begin
    //первый разряд входного числа
    case(f_eight)
        3'o0: value[3:0] = 4'd0;
        3'o1: value[3:0] = 4'd1;
        3'o2: value[3:0] = 4'd2;
        3'o3: value[3:0] = 4'd3;
        3'o4: value[3:0] = 4'd4;
        3'o5: value[3:0] = 4'd5;
        3'o6: value[3:0] = 4'd6;
        3'o7: value[3:0] = 4'd7;
    endcase
    //второй разряд входного числа
    case(s_eignt)
        3'o0: value[7:4] = 4'd0;
        3'o1: value[7:4] = 4'd1;
        3'o2: value[7:4] = 4'd2;
        3'o3: value[7:4] = 4'd3;
        3'o4: value[7:4] = 4'd4;
        3'o5: value[7:4] = 4'd5;
        3'o6: value[7:4] = 4'd6;
        3'o7: value[7:4] = 4'd7;
    endcase
end
endmodule
//На вход подаем значение в двоичном коде. 
//В процессе этого модуля переводим его в ВОСЬМЕРИЧНОЕ представление, смотрим каждый разряд и перебираем все цифры,
//присваивая нужный адрес в chars.v, его всовываем в выделенное место на экране (сделать в ROM отдельно)
//Также для теста сделаю счетчик до 15, значение которого и буду передавать на ROM --> чтобы соблюсти правильность сигналов, реализую счетчик в топе.