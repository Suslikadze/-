`timescale 1ns / 1ps
module char_ROM(
    input clk,
    input en,
    input line,
    input pixels_in,
    output pixels_out,
    output end_of_sumbol,
    output end_of_ROM
);
////////////////////////////////////////////////////////// 

